typedef enum {RED, GREEN, IVORY, YELLOW, BLUE ,} color_e ;

typedef enum {ENGLISH, SPANISH, UKRAINE, NORWAY, JAPANESE} country_e ;

typedef enum {DOG, SNAILS, FOX, HORSE, ZEBRA } pet_e;

typedef enum {COFFEE, TEA, MILK, ORANGE_JUICE, WATER } drink_e ;

typedef enum {OLD_GOLD, KOOL, CHESTERFIELD, LUCKY_STRIKE, PARLIAMENT}  smoke_e;
